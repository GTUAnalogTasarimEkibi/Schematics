** sch_path: /foss/design/xschem (copy)/folded_enes_fd.sch
**.subckt folded_enes_fd VDD VSS MINUS PLUS OUT OUTN
*.iopin VDD
*.iopin VSS
*.iopin MINUS
*.iopin PLUS
*.iopin OUT
*.iopin OUTN
V1 PLUS GND 0.9
V4 MINUS GND 0.9
V5 VSS GND 0
V2 VDD GND 1.8
XM7 net1 net9 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=26 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3
XM8 net2 Vcm1 net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM9 net4 net9 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=26 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3
XM10 net5 Vcm1 net4 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM11 net2 Vcm2 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM12 net3 Vcm3 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM13 net5 Vcm2 net6 VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM14 net6 Vcm3 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM15 net4 MINUS net7 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=30 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM16 net1 PLUS net7 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=30 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM18 net8 net8 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
I1 net9 net8 2.1m
XM19 net9 net9 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM20 OUT net9 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM21 OUT net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=29 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=11 m=11
C1 OUT net3 1.9p m=1
.save  v(out)
.save  v(vcm1)
.save  v(vcm2)
.save  v(net5)
.save  v(net9)
.save  v(net4)
.save  v(net1)
.save  v(net7)
.save  v(net8)
.save  v(net9)
V3 Vcm1 GND 0.3
V6 Vcm2 GND 0.9
.save  v(net6)
.save  v(net3)
XM1 OUTN net5 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=29 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=11 m=11
XM2 OUTN net9 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
C2 OUTN net6 1.9p m=1
V7 Vcm3 GND 0.67191645
.save  v(vcm3)
.save  v(outn)
.save  v(net9)
.save  v(net6)
XM17 net7 net8 VSS GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
.save  v(net2)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control

save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]

save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[gds]

save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[gds]

save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvtv[vdsat]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[gds]

save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm13.msky130_fd_pr__nfet_01v8_lvt[gds]

save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm14.msky130_fd_pr__nfet_01v8_lvt[gds]

save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm15.msky130_fd_pr__nfet_01v8_lvt[gds]

save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm17.msky130_fd_pr__nfet_01v8_lvt[gds]

save @m.xm18.msky130_fd_pr__nfet_01v8[gm]
save @m.xm18.msky130_fd_pr__nfet_01v8[vth]
save @m.xm18.msky130_fd_pr__nfet_01v8[vdsat]
save @m.xm18.msky130_fd_pr__nfet_01v8[vds]
save @m.xm18.msky130_fd_pr__nfet_01v8[id]
save @m.xm18.msky130_fd_pr__nfet_01v8[gds]

save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm19.msky130_fd_pr__pfet_01v8_lvt[gds]

save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[vth]
save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm20.msky130_fd_pr__pfet_01v8_lvt[gds]

save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[vth]
save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm21.msky130_fd_pr__nfet_01v8_lvt[gds]

save all

op
write folded_enes_fd.raw
*.dc Vcm3 Gnd 0.68 0.7 0.002


.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
